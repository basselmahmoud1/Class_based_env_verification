virtual class class_base;
    // `define DEBUG
    protected static event finished_monitoring;
    protected static event finished_driving;
    // protected static event Monitor_now;
    protected static virtual MEM_IF vif_associative [string];
    // protected static class_based_transaction FIFO_trans_handle [$];
endclass